module vga_pic(  
    input wire vga_clk,       // Input working clock, frequency 25MHz  
    input wire sys_rst_n,     // Input reset signal, active low  
    input wire [9:0] pix_x,   // Input pixel X coordinate in the active display area  
    input wire [9:0] pix_y,   // Input pixel Y coordinate in the active display area  

    output reg [15:0] pix_data // Output pixel color information  
);  

    // Parameter definitions  
    parameter CHAR_B_H = 10'd192; // Character start X coordinate  
    parameter CHAR_B_V = 10'd208; // Character start Y coordinate  

    parameter CHAR_W = 10'd256;   // Character width  
    parameter CHAR_H = 10'd64;    // Character height  

    parameter YELLOW = 16'hFFE0;  // Yellow color  
    parameter WHITE = 16'hFFFF;   // White color  
    parameter BLUE = 16'h1C3F;    // Blue color  

    // Internal signal definitions  
    wire [9:0] char_x;            // Character display X coordinate  
    wire [9:0] char_y;            // Character display Y coordinate  

    // Character data storage  
    reg [255:0] char [63:0];      // Character data array  

// Initialize character data   
always@(posedge vga_clk)  
begin  
char [ 0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [ 1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [ 2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [ 3] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [ 4] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [ 5] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [ 6] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [ 7] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [ 8] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [ 9] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [10] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [11] <= 256'h00000000000000000000000000000000000001FFC00000000000000000000000;
char [12] <= 256'h0000FF80000FF8000001FC0001FC000000001FFFFE000000000FFFFFFFF00000;
char [13] <= 256'h0000FF80001FF8000001FC0001FC000000007FFFFF000000000FFFFFFFF00000;
char [14] <= 256'h0000FFC0001FF8000001FC0001FC00000000FFFFFF000000000FFFFFFFF00000;
char [15] <= 256'h0000FFC0003FF8000001FC0001FC00000001FFFFFF000000000FFFFFFFF00000;
char [16] <= 256'h0000FFE0003FF8000001FC0001FC00000003FE0000000000000000FE00000000;
char [17] <= 256'h0000FFE0003FF8000001FC0001FC00000003F80000000000000000FE00000000;
char [18] <= 256'h0000FFF0007FF8000001FC0001FC00000003F80000000000000000FE00000000;
char [19] <= 256'h0001FFF0007DF8000001FC0001FC00000007F00000000000000000FE00000000;
char [20] <= 256'h0001FDF800FDF8000001FC0001FC00000007F00000000000000000FE00000000;
char [21] <= 256'h0001FDF800F9F8000001FC0001FC00000007F00000000000000000FE00000000;
char [22] <= 256'h0001FCFC01F9F8000001FC0001FC00000007F80000000000000000FE00000000;
char [23] <= 256'h0001FCFC01F1F8000001FC0001FC00000003F80000000000000000FE00000000;
char [24] <= 256'h0001FC7C03F1F8000001FC0001FC00000003FC0000000000000000FE00000000;
char [25] <= 256'h0001FC7E03E1FC000001FC0001FC00000003FF8000000000000000FE00000000;
char [26] <= 256'h0001FC3E07E1FC000001FC0001FC00000001FFF000000000000000FE00000000;
char [27] <= 256'h0001FC3F07C1FC000001FC0001FC00000000FFFF00000000000000FE00000000;
char [28] <= 256'h0001F81F0FC1FC000001FC0001FC000000003FFFE0000000000000FE00000000;
char [29] <= 256'h0001F81F8F81FC000001FC0001FC000000000FFFF8000000000000FE00000000;
char [30] <= 256'h0001F80F9F81FC000001FC0001FC0000000001FFFE000000000000FE00000000;
char [31] <= 256'h0001F80FDF01FC000001FC0001FC00000000001FFF000000000000FE00000000;
char [32] <= 256'h0001F807FF01FC000001FC0001FC000000000003FF800000000000FE00000000;
char [33] <= 256'h0001F807FE01FC000001FC0001FC000000000000FF800000000000FE00000000;
char [34] <= 256'h0001F807FE01FC000001FC0001FC0000000000003F800000000000FE00000000;
char [35] <= 256'h0003F803FC01FC000001FC0001FC0000000000003FC00000000000FE00000000;
char [36] <= 256'h0003F803FC01FC000001FC0001FC0000000000001FC00000000000FE00000000;
char [37] <= 256'h0003F801F801FC000001FC0001FC0000000000001FC00000000000FE00000000;
char [38] <= 256'h0003F8000001FC000001FC0003FC0000000000001FC00000000000FE00000000;
char [39] <= 256'h0003F8000001FC000001FC0003F80000000000003FC00000000000FE00000000;
char [40] <= 256'h0003F8000001FC000001FE0007F80000000000003F800000000000FE00000000;
char [41] <= 256'h0003F8000001FC000000FF000FF00000000000007F800000000000FE00000000;
char [42] <= 256'h0003F8000001FC000000FFC03FF0000000038003FF000000000000FE00000000;
char [43] <= 256'h0003F8000001FC0000007FFFFFE000000003FFFFFF000000000000FE00000000;
char [44] <= 256'h0003F8000001FC0000003FFFFFC000000003FFFFFE000000000000FE00000000;
char [45] <= 256'h0003F8000001FC0000000FFFFF8000000003FFFFF8000000000000FE00000000;
char [46] <= 256'h0003F8000000FC00000003FFFC0000000001FFFFE0000000000000FE00000000;
char [47] <= 256'h00000000000000000000000700000000000000F0000000000000000000000000;
char [48] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [49] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [50] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [51] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [52] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [53] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [54] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [55] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [56] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [57] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [58] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [59] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [60] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char [63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
end  

 // Calculate character display coordinates  
    assign char_x = (pix_x >= CHAR_B_H && pix_x < (CHAR_B_H + CHAR_W)) ? (pix_x - CHAR_B_H) : 10'h3FF;  
    assign char_y = (pix_y >= CHAR_B_V && pix_y < (CHAR_B_V + CHAR_H)) ? (pix_y - CHAR_B_V) : 10'h3FF;  

    // Determine pixel color based on character data  
    always @(posedge vga_clk or negedge sys_rst_n) begin  
        if (!sys_rst_n) begin  
            pix_data <= YELLOW; // Default color on reset  
        end else if (char_x != 10'h3FF && char_y != 10'h3FF && char[char_y][255 - char_x]) begin  
            pix_data <= BLUE;   // Display blue if character pixel is set  
        end else begin  
            pix_data <= YELLOW; // Display yellow otherwise  
        end  
    end  

endmodule  
